*/////////////////////////////////////////////////////
* LTC7652  Chopper-Stabilised Operational Amplifier //
*/////////////////////////////////////////////////////
*
* connections:     non-inverting input
*                  |   inverting input
*                  |   |   positive power supply
*                  |   |   |   negative power supply
*                  |   |   |   |   output
*                  |   |   |   |   |
*                  |   |   |   |   |
.SUBCKT LTC7652    3   2   7   4   6 
X_LTC7652 3 2 7 4 6 LTC1052
.ENDS LTC7652
*
***
*
.SUBCKT LTC1052    3 2 7 4 6 
* INPUT
IB1 2 7 -10P
IB2 3 7 10P
RD1 4 80 4.4210E+03
RD2 4 90 4.4210E+03
M1 80 2 12 12 PM1 
M2 90 3 12 12 PM2 
CIN 2 3 5.0000E-12
DG1 2 7 DMG1
DG2 3 7 DMG2
C1 80 90 1.5000E-11
ISS 7 12 1.2000E-04
CS 12 0 7.5000E-12
* INTERMEDIATE 
GCM 0 8 12 0 2.2619E-11
GA 8 0 80 90 2.2619E-04
R2 8 0 1.0000E+05
C2 1 8 3.0000E-11
GB 1 0 8 0 7.0253E+03
RO2 1 0 1.9900E+02
* OUTPUT 
RSO 1 6 1.0000E+00
ECL 18 0 1 6 1.7955E+02
GCL 0 8 20 0 1.0000E+00
RCL 20 0 1.0000E+01
D1 18 19 DM1 
VOD1 19 20 0.0000E+00
D2 20 21 DM1 
VOD2 21 18 1.7955E+00
* 
D3A 131 70 DM3 
D3B 13 131 DM3 
GPL 0 8 70 7 1.0000E+00
VC 13 6 1.4332E+00
RPLA 7 70 1.0000E+01
RPLB 7 131 1.0000E+03
D4A 60 141 DM3 
D4B 141 14 DM3 
GNL 0 8 60 4 1.0000E+00
VE 6 14 1.4332E+00
RNLA 60 4 1.0000E+01
RNLB 141 4 1.0000E+03
* 
IP 7 4 1.5800E-03
DSUB 4 7 DM2 
* MODELS 
.MODEL PM1 PMOS (KP=4.2637E-04 VTO=-1.1000000E+00)
.MODEL PM2 PMOS (KP=4.2637E-04 VTO=-1.1000005E+00)
.MODEL DM1 D (IS=1.0000E-20)
.MODEL DM2 D (IS=8.0000E-16 BV=1.9800E+01)
.MODEL DM3 D (IS=1.0000E-16)
.MODEL DMG1 D (IS=7E-12 N=2.31)
.MODEL DMG2 D (IS=6.3E-12 N=2.31)
.ENDS LTC1052